library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

use work.ctrl_common.all;

entity bofp1 is
    generic (
        G_CFG_WIDTH: integer := 12; -- Width of config entries,
        G_ADC_WIDTH: integer := 16 -- Width/resoluton of ADC readouts
    );
    port (
        i_clk: in std_logic;

        o_ccd_sh: out std_logic;
        o_ccd_mclk: out std_logic;
        o_ccd_icg: out std_logic;
        o_ccd_busy: out std_logic;

        i_adc_eoc: in std_logic;
        o_adc_stconv: out std_logic;

        o_fifo_wmark: out std_logic;

        i_spi_main_miso: in std_logic;
        o_spi_main_mosi: out std_logic;
        o_spi_main_sclk: out std_logic;
        o_spi_main_cs_n: out std_logic;

        i_spi_sub_sclk: in std_logic;
        i_spi_sub_cs_n: in std_logic;
        i_spi_sub_mosi: in std_logic;
        o_spi_sub_miso: out std_logic
    );
end entity bofp1;

architecture structural of bofp1 is
    signal r_clk_main: std_logic;

    signal r_rst: std_logic;
    signal r_rst_n: std_logic;
    signal r_rst_en: std_logic;

    signal r_ccd_start: std_logic; -- Passed to control module
    signal r_ccd_data_rdy: std_logic;

    signal r_adc_spi_sclk: std_logic;
    signal r_adc_spi_data: std_logic_vector(G_ADC_WIDTH-1 downto 0);
    signal r_adc_spi_rdy: std_logic; -- Ready to read out

    signal r_ctrl_fifo_rd_en: std_logic;
    signal r_ctrl_fifo_val: std_logic_vector(G_ADC_WIDTH-1 downto 0);

    signal r_fifo_empty: std_logic;

    signal r_regmap: t_regmap;

    -- FIFO generated by Vivado, used for storing the raw voltages from
    -- the CCD ADC.
    -- 1024x16, full, empty flag
    -- Independent clock distributed RAM
    component fifo_data is
        port (
            rst: in std_logic;
            wr_clk: in std_logic;
            rd_clk: in std_logic;
            din: in std_logic_vector(G_ADC_WIDTH-1 downto 0);
            wr_en: in std_logic;
            rd_en: in std_logic;
            dout: out std_logic_vector(G_ADC_WIDTH-1 downto 0);
            full: out std_logic;
            empty: out std_logic;
            prog_full: out std_logic
        );
    end component fifo_data;

    -- Clocking wizard generated by Vivado
    -- clk_in1: 100 MHz
    -- sclk_adc: SCLK for the SPI interaction with the ADC. 25MHz
    component clk_wizard is
        port (
            clk_in1: in std_logic;
            main: out std_logic;
            sclk_adc: out std_logic;
            locked: out std_logic
        );
    end component clk_wizard;
begin
    r_rst_n <= not r_rst;
    o_spi_main_sclk <= r_adc_spi_sclk;

    u_reset: entity work.reset(rtl)
        generic map(
            G_CYC_COUNT => 4
        )
        port map(
            i_clk => i_clk,
            i_en => r_rst_en,
            o_rst => r_rst
        );

    u_clk: clk_wizard
        port map(
            clk_in1 => i_clk,
            main => r_clk_main,
            sclk_adc => r_adc_spi_sclk
        );

    u_ccd: entity work.tcd1304(rtl) generic map(
        G_CLK_FREQ => 100_000_000 -- TODO
    )
    port map(
        i_clk => r_clk_main,
        i_rst_n => r_rst_n,
        i_start => r_ccd_start,
        i_psc_div => r_regmap.clkdiv(7 downto 3), 
        i_sh_div => r_regmap.shdiv,
        i_mclk_div => r_regmap.clkdiv(2 downto 0),

        o_pin_sh => o_ccd_sh,
        o_pin_mclk => o_ccd_mclk,
        o_pin_icg => o_ccd_icg,
        o_data_rdy => r_ccd_data_rdy,
        o_ccd_busy => o_ccd_busy
    );

    u_adc: entity work.ads8329(rtl) port map(
        i_clk => r_clk_main,
        i_rst_n => r_rst_n,
        i_start => r_ccd_data_rdy,

        i_pin_eoc => i_adc_eoc,
        o_pin_stconv => o_adc_stconv,

        i_miso => i_spi_main_miso,
        i_sclk => r_adc_spi_sclk,
        o_mosi => o_spi_main_mosi,
        o_cs_n => o_spi_main_cs_n,

        o_data => r_adc_spi_data,
        o_rdy => r_adc_spi_rdy
    );

    u_fifo_data: fifo_data port map (
        rst => r_rst,
        wr_clk => r_clk_main,
        rd_clk => i_spi_sub_sclk,
        wr_en => r_adc_spi_rdy,
        din => r_adc_spi_data,
        rd_en => r_ctrl_fifo_rd_en,
        dout => r_ctrl_fifo_val,
        empty => r_fifo_empty,
        prog_full => o_fifo_wmark
    );

    u_ctrl: entity work.ctrl(behaviour) port map(
        i_clk => r_clk_main,
        i_rst_n => r_rst_n,
        o_ccd_sample => r_ccd_start,
        o_rst => r_rst_en,

        i_sclk => i_spi_sub_sclk,
        i_cs_n => i_spi_sub_cs_n,
        i_mosi => i_spi_sub_mosi,
        o_miso => o_spi_sub_miso,

        i_fifo_empty => r_fifo_empty,
        i_fifo_data => r_ctrl_fifo_val,
        o_fifo_rd => r_ctrl_fifo_rd_en,

        o_regmap => r_regmap
    );

end architecture structural;
