library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity bofp1 is
    generic (
        G_CFG_WIDTH: integer := 12; -- Width of config entries,
        G_ADC_WIDTH: integer := 16; -- Width/resoluton of ADC readouts
        G_CTRL_WIDTH: integer := 16 -- Width of ctrl codes
    );
    port (
        i_clk: in std_logic;
        i_rst: in std_logic;

        o_ccd_sh: out std_logic;
        o_ccd_mclk: out std_logic;
        o_ccd_icg: out std_logic;

        i_adc_eoc: in std_logic;
        o_adc_stconv: out std_logic;

        i_spi_main_miso: in std_logic;
        o_spi_main_mosi: out std_logic;
        o_spi_main_sclk: out std_logic;

        i_spi_sub_sclk: in std_logic;
        i_spi_sub_cs_n: in std_logic;
        i_spi_sub_mosi: in std_logic;
        o_spi_sub_miso: out std_logic
    );
end entity bofp1;

architecture structural of bofp1 is
    signal r_rst_n: std_logic;

    signal r_ccd_start: std_logic; -- Passed to control module
    signal r_ccd_data_rdy: std_logic;

    signal r_adc_spi_en: std_logic; -- Start read
    signal r_adc_spi_data: std_logic_vector(G_ADC_WIDTH-1 downto 0);
    signal r_adc_spi_rdy: std_logic; -- Ready to read out

    signal r_ctrl_wr_en: std_logic;
    signal r_ctrl_wr_data: std_logic_vector(G_CTRL_WIDTH-1 downto 0);
    signal r_ctrl_rd_en: std_logic;
    signal r_ctrl_rd_data: std_logic_vector(G_CTRL_WIDTH-1 downto 0);
    signal r_ctrl_fifo_rd_en: std_logic;
    signal r_ctrl_fifo_val: std_logic_vector(G_ADC_WIDTH-1 downto 0);

    signal r_spi_sub_rdy: std_logic;
    signal r_spi_sub_data_rd: std_logic_vector(G_CTRL_WIDTH-1 downto 0);
    signal r_spi_sub_data_wr: std_logic_vector(G_CTRL_WIDTH-1 downto 0);

    -- FIFO generated by Vivado, used for storing the raw voltages from
    -- the CCD ADC.
    -- 1024x16, full, empty flag
    -- Independent clock distributed RAM
    component fifo_generator_0 is
        port (
            rst: in std_logic;
            wr_clk: in std_logic;
            rd_clk: in std_logic;
            din: in std_logic_vector(G_ADC_WIDTH-1 downto 0);
            wr_en: in std_logic;
            rd_en: in std_logic;
            dout: out std_logic_vector(G_ADC_WIDTH-1 downto 0);
            full: out std_logic;
            empty: out std_logic
        );
    end component fifo_generator_0;

    -- FIFO generated by Vivado, used for crossing the configuration
    -- parameters from the SCLK domain to the CLK domain.
    -- 16x16, full, empty flag
    -- Independet clock distributed RAM
    component fifo_ctrl is
        port (
            rst: in std_logic;
            wr_clk: in std_logic;
            rd_clk: in std_logic;
            din: in std_logic_vector(G_CTRL_WIDTH-1 downto 0);
            wr_en: in std_logic;
            rd_en: in std_logic;
            dout: out std_logic_vector(G_CTRL_WIDTH-1 downto 0);
            full: out std_logic;
            empty: out std_logic
        );
    end component fifo_ctrl;
begin
    r_rst_n <= not i_rst;

    u_ccd: entity work.tcd1304(rtl) generic map(
        G_CFG_WIDTH => G_CFG_WIDTH,
        G_CLK_FREQ => 100_000_000 -- TODO
    )
    port map(
        i_clk => i_clk,
        i_rst_n => r_rst_n,
        i_start => r_ccd_start,
        i_sh_div => std_logic_vector(to_unsigned(50, G_CFG_WIDTH)), -- TODO
        i_mclk_div => std_logic_vector(to_unsigned(50, G_CFG_WIDTH)), -- TODO

        o_pin_sh => o_ccd_sh,
        o_pin_mclk => o_ccd_mclk,
        o_pin_icg => o_ccd_icg,
        o_data_rdy => r_ccd_data_rdy
    );

    u_adc: entity work.ads8329(rtl) generic map(
        G_CLK_DIV => 10
    )
    port map(
        i_clk => i_clk,
        i_rst_n => r_rst_n,
        i_start => r_ccd_data_rdy,

        i_pin_eoc => i_adc_eoc,
        o_pin_stconv => o_adc_stconv,

        o_rd_en => r_adc_spi_en
    );

    u_adc_spi: entity work.spi_main(rtl) generic map(
        G_DATA_WIDTH => G_ADC_WIDTH,
        G_CLK_DIV => 4
    )
    port map(
        i_clk => i_clk,
        i_rst_n => r_rst_n,
        i_rd_en => r_adc_spi_en,
        i_data => "1101000000000000",

        i_miso => i_spi_main_miso,
        o_mosi => o_spi_main_mosi,
        o_sclk => o_spi_main_sclk,

        o_data => r_adc_spi_data,
        o_rd_en => r_adc_spi_rdy
    );

    u_fifo_data: fifo_generator_0 port map (
        rst => i_rst,
        wr_clk => i_clk,
        rd_clk => i_spi_sub_sclk,
        wr_en => r_adc_spi_rdy,
        din => r_adc_spi_data,
        rd_en => r_ctrl_fifo_rd_en,
        dout => r_ctrl_fifo_val
    );

    u_ctrl_spi: entity work.spi_sub(rtl) generic map(
        G_DATA_WIDTH => G_CTRL_WIDTH
    )
    port map(
        i_sclk => i_spi_sub_sclk,
        i_arst_n => r_rst_n,
        i_data => r_spi_sub_data_wr,
        
        i_mosi => i_spi_sub_mosi,
        i_cs_n => i_spi_sub_cs_n,
        o_miso => o_spi_sub_miso,

        o_data => r_spi_sub_data_rd,
        o_rdy => r_spi_sub_rdy
    );

    /*
    ctrl port map(
        i_clk
        i_rst

        i_spi_sub_data_rd

        o => r_ctrl_wr_en
        o => r_ctrl_wr_data

        i => r_ctrl_rd_en
        i => r_ctrl_rd_data


        o_spi_sub_data_wr
    )
    */

    u_fifo_ctrl: fifo_ctrl port map(
        rst => i_rst,
        wr_clk => i_spi_sub_sclk,
        rd_clk => i_clk,
        wr_en => r_ctrl_wr_en,
        din => r_ctrl_wr_data,
        rd_en => r_ctrl_rd_en,
        dout => r_ctrl_rd_data
    );

end architecture structural;
